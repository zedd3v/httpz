module httpz

pub fn test() string {
	return 'hello'
}
